`timescale 1ns/1ps

module EVP_FSM_3 
		#(parameter buffer_size = 1024)(
		input clk, rst,
		input rst_instr,
		input start_evp,
		input [2 : 0] A,
		input [15 : 0] x,
		input [15 : 0] c_i,
		input [4 : 0] N,
		input [log2(buffer_size)-1 : 0] rd_addr_data, 
		output reg en_rd_data,
		output reg en_rd_S,
		output reg en_rd_N,
		output reg [log2(buffer_size)-1 : 0] rd_addr_data_updated,
		output [6 : 0] rd_addr_S,
		output reg [2 : 0] rd_addr_N,
		output reg done_evp,
		output reg [31 : 0] result,
		output reg [31 : 0] status);

		reg [2 : 0] state, next_state;
		reg [31 : 0] next_result;
		reg [31 : 0] next_status;
		reg [3 : 0] S_idx_counter, next_S_idx_counter;
		reg [3 : 0] exp_counter, next_exp_counter;
		reg [31 : 0] monomial, next_monomial;
		reg [31 : 0] sum, next_sum;
		reg [log2(buffer_size)-1 : 0] next_rd_addr_data;

	localparam STATE_START = 3'b000, STATE_COMPUTE0 = 3'b001, 
				STATE_COMPUTE1 = 3'b010, STATE_COMPUTE2 = 3'b011,
				STATE_ERROR = 3'b100, STATE_END = 3'b101;

assign rd_addr_data = rd_addr_data_updated;
assign rd_addr_S = A * 11 + S_idx_counter;

	always @(posedge clk, negedge rst)
		if (! rst || ! rst_instr) begin
			$display("rst");
			state <= STATE_START;
			monomial <= 1;
			sum <= 0;
			S_idx_counter <= 0;
			exp_counter <= 0;
			rd_addr_data_updated <= 0;
			result <= 0;
			status <= 32'b11111111111111111111111111111111;
		end
		else begin
			$display("state = ", state, ", next_state = ", next_state);
			state <= next_state;
			monomial <= next_monomial;
			sum <= next_sum;
			S_idx_counter <= next_S_idx_counter;
			exp_counter <= next_exp_counter;
			rd_addr_data_updated <= next_rd_addr_data;
			result <= next_result;
			status <= next_status;
		end

	always @(state, start_evp, S_idx_counter, N)
		case (state)
			STATE_START:
			begin
				if (start_evp)
					next_state <= STATE_COMPUTE0;
				else
					next_state <= STATE_START;
			end

			STATE_COMPUTE0:
				if (N == 5'b11111)
					next_state <= STATE_ERROR;
				else
					next_state <= STATE_COMPUTE1;

			STATE_COMPUTE1:
			begin
				if (S_idx_counter > N) begin
					$display("S_idx_counter > N: ", S_idx_counter, " > ", N);
					next_state <= STATE_END;
				end
				else if (exp_counter == S_idx_counter) begin
					$display("hit condition exp_counter == S_idx_counter");
					next_state <= STATE_COMPUTE2;
				end
				else begin
					$display("exp_counter = ", exp_counter, ", S_idx_counter = ", S_idx_counter);
					next_state <= STATE_COMPUTE1;
				end
			end

			STATE_COMPUTE2:
			begin
				//if (S_idx_counter > N)
				//	next_state <= STATE_END;
				//else
				next_state <= STATE_COMPUTE1;
			end

			STATE_ERROR:
				next_state <= STATE_END;

			STATE_END:
				next_state <= STATE_START;
	
		endcase

	always @(state, start_evp, rd_addr_data, rd_addr_data_updated, 
				S_idx_counter, exp_counter, c_i, x, monomial, sum, result, 
				status)
		case (state)
			STATE_START:
			begin
				done_evp <= 0;
				en_rd_data <= 0;
				en_rd_S <= 0;
				en_rd_N <= 0;
				next_monomial <= 1;
				next_sum <= 0;
				next_S_idx_counter <= 0;
				next_exp_counter <= 0;
				next_rd_addr_data <= rd_addr_data;
				rd_addr_N <= rd_addr_N;
				next_result <= 0;
				next_status <= 32'b11111111111111111111111111111111;
			end

			STATE_COMPUTE0:
			begin
				done_evp <= 0;
				en_rd_data <= 1;
				en_rd_S <= 1;
				en_rd_N <= 1;
				next_monomial <= 1;
				next_sum <= sum;
				next_S_idx_counter <= S_idx_counter;
				next_exp_counter <= exp_counter;
				next_rd_addr_data <= rd_addr_data_updated + 1;
				rd_addr_N <= A;
				next_result <= result;
				next_status <= status;
			end

			STATE_COMPUTE1:
			begin
				done_evp <= 0;
				en_rd_data <= 0;
				en_rd_S <= 0;
				en_rd_N <= 0;
				next_monomial <= monomial * x;
				next_sum <= sum;
				next_S_idx_counter <= S_idx_counter;
				$display("S_idx_counter = ", S_idx_counter, ", next_S_idx_counter = ", next_S_idx_counter);
				next_exp_counter <= exp_counter + 1;
				$display("exp_counter = ", exp_counter, ", next_exp_counter = ", next_exp_counter);
				next_rd_addr_data <= rd_addr_data_updated;
				rd_addr_N <= rd_addr_N;
				next_result <= result;
				next_status <= status; 
			end

			STATE_COMPUTE2:
			begin
				done_evp <= 0;
				en_rd_data <= 0;
				en_rd_S <= 1;
				en_rd_N <= 0;
				next_monomial <= 1;
				next_sum <= sum + monomial * c_i;
				next_S_idx_counter <= S_idx_counter + 1;
				$display("S_idx_counter = ", S_idx_counter, ", next_S_idx_counter = ", next_S_idx_counter);
				next_exp_counter <= 0;
				$display("exp_counter = ", exp_counter, ", next_exp_counter = ", next_exp_counter);
				next_rd_addr_data <= rd_addr_data_updated;
				rd_addr_N <= rd_addr_N;
				next_result <= result;
				next_status <= status;
			end

			STATE_ERROR:
			begin
				done_evp <= 0;
				en_rd_data <= 0;
				en_rd_S <= 0;
				en_rd_N <= 0;
				next_monomial <= monomial;
				next_sum <= sum;
				next_S_idx_counter <= S_idx_counter;
				next_exp_counter <= exp_counter;
				next_rd_addr_data <= rd_addr_data_updated;
				rd_addr_N <= rd_addr_N;
				next_result <= 0;
				next_status <= 2'b10;
			end

			STATE_END:
			begin
				done_evp <= 1;
				en_rd_data <= 0;
				en_rd_S <= 0;
				en_rd_N <= 0;
				next_monomial <= monomial;
				next_sum <= sum;
				next_S_idx_counter <= S_idx_counter;
				next_exp_counter <= exp_counter;
				next_rd_addr_data <= rd_addr_data_updated;
				rd_addr_N <= rd_addr_N;
				next_result <= sum;
				next_status <= 0;
			end
		endcase

	function integer log2;
    input [31 : 0] value;
     integer i;
    begin
          if(value==1)
                log2=1;
          else
              begin
              i = value - 1;
              for (log2 = 0; i > 0; log2 = log2 + 1) begin
                    i = i >> 1;
              end
              end
    end
    endfunction

endmodule	
